// Output module generated using c++
// sends final state-vector to arduino
module output_2qb #(
parameter N = 16
)
(
input [N-1:0] psi_f [0:287],
input wire i_clock,
input wire listener_flag,
output wire[7:0] out,
output wire parity
);

// used for iterating through output
integer n_num = 576;
integer i_num = 0;
reg [7:0] out_reg; // for assigning numbers in always block
assign out[7:0] = out_reg[7:0];
reg parity_reg;
assign parity = parity_reg;

// intialization of values
initial begin
    out_reg <= 8'b10001011;
    parity_reg <= 1'b0;
end


// transfer data to arduino
always @ (posedge listener_flag)
begin
    case(i_num)
    0: begin
         out_reg[7:0] <= psi_f[0][15:8];
         parity_reg <= ^psi_f[0][15:8];
       end
    1: begin
         out_reg[7:0] <= psi_f[0][7:0];
         parity_reg <= ^psi_f[0][7:0];
       end
    2: begin
         out_reg[7:0] <= psi_f[1][15:8];
         parity_reg <= ^psi_f[1][15:8];
       end
    3: begin
         out_reg[7:0] <= psi_f[1][7:0];
         parity_reg <= ^psi_f[1][7:0];
       end
    4: begin
         out_reg[7:0] <= psi_f[2][15:8];
         parity_reg <= ^psi_f[2][15:8];
       end
    5: begin
         out_reg[7:0] <= psi_f[2][7:0];
         parity_reg <= ^psi_f[2][7:0];
       end
    6: begin
         out_reg[7:0] <= psi_f[3][15:8];
         parity_reg <= ^psi_f[3][15:8];
       end
    7: begin
         out_reg[7:0] <= psi_f[3][7:0];
         parity_reg <= ^psi_f[3][7:0];
       end
    8: begin
         out_reg[7:0] <= psi_f[4][15:8];
         parity_reg <= ^psi_f[4][15:8];
       end
    9: begin
         out_reg[7:0] <= psi_f[4][7:0];
         parity_reg <= ^psi_f[4][7:0];
       end
    10: begin
         out_reg[7:0] <= psi_f[5][15:8];
         parity_reg <= ^psi_f[5][15:8];
       end
    11: begin
         out_reg[7:0] <= psi_f[5][7:0];
         parity_reg <= ^psi_f[5][7:0];
       end
    12: begin
         out_reg[7:0] <= psi_f[6][15:8];
         parity_reg <= ^psi_f[6][15:8];
       end
    13: begin
         out_reg[7:0] <= psi_f[6][7:0];
         parity_reg <= ^psi_f[6][7:0];
       end
    14: begin
         out_reg[7:0] <= psi_f[7][15:8];
         parity_reg <= ^psi_f[7][15:8];
       end
    15: begin
         out_reg[7:0] <= psi_f[7][7:0];
         parity_reg <= ^psi_f[7][7:0];
       end
    16: begin
         out_reg[7:0] <= psi_f[8][15:8];
         parity_reg <= ^psi_f[8][15:8];
       end
    17: begin
         out_reg[7:0] <= psi_f[8][7:0];
         parity_reg <= ^psi_f[8][7:0];
       end
    18: begin
         out_reg[7:0] <= psi_f[9][15:8];
         parity_reg <= ^psi_f[9][15:8];
       end
    19: begin
         out_reg[7:0] <= psi_f[9][7:0];
         parity_reg <= ^psi_f[9][7:0];
       end
    20: begin
         out_reg[7:0] <= psi_f[10][15:8];
         parity_reg <= ^psi_f[10][15:8];
       end
    21: begin
         out_reg[7:0] <= psi_f[10][7:0];
         parity_reg <= ^psi_f[10][7:0];
       end
    22: begin
         out_reg[7:0] <= psi_f[11][15:8];
         parity_reg <= ^psi_f[11][15:8];
       end
    23: begin
         out_reg[7:0] <= psi_f[11][7:0];
         parity_reg <= ^psi_f[11][7:0];
       end
    24: begin
         out_reg[7:0] <= psi_f[12][15:8];
         parity_reg <= ^psi_f[12][15:8];
       end
    25: begin
         out_reg[7:0] <= psi_f[12][7:0];
         parity_reg <= ^psi_f[12][7:0];
       end
    26: begin
         out_reg[7:0] <= psi_f[13][15:8];
         parity_reg <= ^psi_f[13][15:8];
       end
    27: begin
         out_reg[7:0] <= psi_f[13][7:0];
         parity_reg <= ^psi_f[13][7:0];
       end
    28: begin
         out_reg[7:0] <= psi_f[14][15:8];
         parity_reg <= ^psi_f[14][15:8];
       end
    29: begin
         out_reg[7:0] <= psi_f[14][7:0];
         parity_reg <= ^psi_f[14][7:0];
       end
    30: begin
         out_reg[7:0] <= psi_f[15][15:8];
         parity_reg <= ^psi_f[15][15:8];
       end
    31: begin
         out_reg[7:0] <= psi_f[15][7:0];
         parity_reg <= ^psi_f[15][7:0];
       end
    32: begin
         out_reg[7:0] <= psi_f[16][15:8];
         parity_reg <= ^psi_f[16][15:8];
       end
    33: begin
         out_reg[7:0] <= psi_f[16][7:0];
         parity_reg <= ^psi_f[16][7:0];
       end
    34: begin
         out_reg[7:0] <= psi_f[17][15:8];
         parity_reg <= ^psi_f[17][15:8];
       end
    35: begin
         out_reg[7:0] <= psi_f[17][7:0];
         parity_reg <= ^psi_f[17][7:0];
       end
    36: begin
         out_reg[7:0] <= psi_f[18][15:8];
         parity_reg <= ^psi_f[18][15:8];
       end
    37: begin
         out_reg[7:0] <= psi_f[18][7:0];
         parity_reg <= ^psi_f[18][7:0];
       end
    38: begin
         out_reg[7:0] <= psi_f[19][15:8];
         parity_reg <= ^psi_f[19][15:8];
       end
    39: begin
         out_reg[7:0] <= psi_f[19][7:0];
         parity_reg <= ^psi_f[19][7:0];
       end
    40: begin
         out_reg[7:0] <= psi_f[20][15:8];
         parity_reg <= ^psi_f[20][15:8];
       end
    41: begin
         out_reg[7:0] <= psi_f[20][7:0];
         parity_reg <= ^psi_f[20][7:0];
       end
    42: begin
         out_reg[7:0] <= psi_f[21][15:8];
         parity_reg <= ^psi_f[21][15:8];
       end
    43: begin
         out_reg[7:0] <= psi_f[21][7:0];
         parity_reg <= ^psi_f[21][7:0];
       end
    44: begin
         out_reg[7:0] <= psi_f[22][15:8];
         parity_reg <= ^psi_f[22][15:8];
       end
    45: begin
         out_reg[7:0] <= psi_f[22][7:0];
         parity_reg <= ^psi_f[22][7:0];
       end
    46: begin
         out_reg[7:0] <= psi_f[23][15:8];
         parity_reg <= ^psi_f[23][15:8];
       end
    47: begin
         out_reg[7:0] <= psi_f[23][7:0];
         parity_reg <= ^psi_f[23][7:0];
       end
    48: begin
         out_reg[7:0] <= psi_f[24][15:8];
         parity_reg <= ^psi_f[24][15:8];
       end
    49: begin
         out_reg[7:0] <= psi_f[24][7:0];
         parity_reg <= ^psi_f[24][7:0];
       end
    50: begin
         out_reg[7:0] <= psi_f[25][15:8];
         parity_reg <= ^psi_f[25][15:8];
       end
    51: begin
         out_reg[7:0] <= psi_f[25][7:0];
         parity_reg <= ^psi_f[25][7:0];
       end
    52: begin
         out_reg[7:0] <= psi_f[26][15:8];
         parity_reg <= ^psi_f[26][15:8];
       end
    53: begin
         out_reg[7:0] <= psi_f[26][7:0];
         parity_reg <= ^psi_f[26][7:0];
       end
    54: begin
         out_reg[7:0] <= psi_f[27][15:8];
         parity_reg <= ^psi_f[27][15:8];
       end
    55: begin
         out_reg[7:0] <= psi_f[27][7:0];
         parity_reg <= ^psi_f[27][7:0];
       end
    56: begin
         out_reg[7:0] <= psi_f[28][15:8];
         parity_reg <= ^psi_f[28][15:8];
       end
    57: begin
         out_reg[7:0] <= psi_f[28][7:0];
         parity_reg <= ^psi_f[28][7:0];
       end
    58: begin
         out_reg[7:0] <= psi_f[29][15:8];
         parity_reg <= ^psi_f[29][15:8];
       end
    59: begin
         out_reg[7:0] <= psi_f[29][7:0];
         parity_reg <= ^psi_f[29][7:0];
       end
    60: begin
         out_reg[7:0] <= psi_f[30][15:8];
         parity_reg <= ^psi_f[30][15:8];
       end
    61: begin
         out_reg[7:0] <= psi_f[30][7:0];
         parity_reg <= ^psi_f[30][7:0];
       end
    62: begin
         out_reg[7:0] <= psi_f[31][15:8];
         parity_reg <= ^psi_f[31][15:8];
       end
    63: begin
         out_reg[7:0] <= psi_f[31][7:0];
         parity_reg <= ^psi_f[31][7:0];
       end
    64: begin
         out_reg[7:0] <= psi_f[32][15:8];
         parity_reg <= ^psi_f[32][15:8];
       end
    65: begin
         out_reg[7:0] <= psi_f[32][7:0];
         parity_reg <= ^psi_f[32][7:0];
       end
    66: begin
         out_reg[7:0] <= psi_f[33][15:8];
         parity_reg <= ^psi_f[33][15:8];
       end
    67: begin
         out_reg[7:0] <= psi_f[33][7:0];
         parity_reg <= ^psi_f[33][7:0];
       end
    68: begin
         out_reg[7:0] <= psi_f[34][15:8];
         parity_reg <= ^psi_f[34][15:8];
       end
    69: begin
         out_reg[7:0] <= psi_f[34][7:0];
         parity_reg <= ^psi_f[34][7:0];
       end
    70: begin
         out_reg[7:0] <= psi_f[35][15:8];
         parity_reg <= ^psi_f[35][15:8];
       end
    71: begin
         out_reg[7:0] <= psi_f[35][7:0];
         parity_reg <= ^psi_f[35][7:0];
       end
    72: begin
         out_reg[7:0] <= psi_f[36][15:8];
         parity_reg <= ^psi_f[36][15:8];
       end
    73: begin
         out_reg[7:0] <= psi_f[36][7:0];
         parity_reg <= ^psi_f[36][7:0];
       end
    74: begin
         out_reg[7:0] <= psi_f[37][15:8];
         parity_reg <= ^psi_f[37][15:8];
       end
    75: begin
         out_reg[7:0] <= psi_f[37][7:0];
         parity_reg <= ^psi_f[37][7:0];
       end
    76: begin
         out_reg[7:0] <= psi_f[38][15:8];
         parity_reg <= ^psi_f[38][15:8];
       end
    77: begin
         out_reg[7:0] <= psi_f[38][7:0];
         parity_reg <= ^psi_f[38][7:0];
       end
    78: begin
         out_reg[7:0] <= psi_f[39][15:8];
         parity_reg <= ^psi_f[39][15:8];
       end
    79: begin
         out_reg[7:0] <= psi_f[39][7:0];
         parity_reg <= ^psi_f[39][7:0];
       end
    80: begin
         out_reg[7:0] <= psi_f[40][15:8];
         parity_reg <= ^psi_f[40][15:8];
       end
    81: begin
         out_reg[7:0] <= psi_f[40][7:0];
         parity_reg <= ^psi_f[40][7:0];
       end
    82: begin
         out_reg[7:0] <= psi_f[41][15:8];
         parity_reg <= ^psi_f[41][15:8];
       end
    83: begin
         out_reg[7:0] <= psi_f[41][7:0];
         parity_reg <= ^psi_f[41][7:0];
       end
    84: begin
         out_reg[7:0] <= psi_f[42][15:8];
         parity_reg <= ^psi_f[42][15:8];
       end
    85: begin
         out_reg[7:0] <= psi_f[42][7:0];
         parity_reg <= ^psi_f[42][7:0];
       end
    86: begin
         out_reg[7:0] <= psi_f[43][15:8];
         parity_reg <= ^psi_f[43][15:8];
       end
    87: begin
         out_reg[7:0] <= psi_f[43][7:0];
         parity_reg <= ^psi_f[43][7:0];
       end
    88: begin
         out_reg[7:0] <= psi_f[44][15:8];
         parity_reg <= ^psi_f[44][15:8];
       end
    89: begin
         out_reg[7:0] <= psi_f[44][7:0];
         parity_reg <= ^psi_f[44][7:0];
       end
    90: begin
         out_reg[7:0] <= psi_f[45][15:8];
         parity_reg <= ^psi_f[45][15:8];
       end
    91: begin
         out_reg[7:0] <= psi_f[45][7:0];
         parity_reg <= ^psi_f[45][7:0];
       end
    92: begin
         out_reg[7:0] <= psi_f[46][15:8];
         parity_reg <= ^psi_f[46][15:8];
       end
    93: begin
         out_reg[7:0] <= psi_f[46][7:0];
         parity_reg <= ^psi_f[46][7:0];
       end
    94: begin
         out_reg[7:0] <= psi_f[47][15:8];
         parity_reg <= ^psi_f[47][15:8];
       end
    95: begin
         out_reg[7:0] <= psi_f[47][7:0];
         parity_reg <= ^psi_f[47][7:0];
       end
    96: begin
         out_reg[7:0] <= psi_f[48][15:8];
         parity_reg <= ^psi_f[48][15:8];
       end
    97: begin
         out_reg[7:0] <= psi_f[48][7:0];
         parity_reg <= ^psi_f[48][7:0];
       end
    98: begin
         out_reg[7:0] <= psi_f[49][15:8];
         parity_reg <= ^psi_f[49][15:8];
       end
    99: begin
         out_reg[7:0] <= psi_f[49][7:0];
         parity_reg <= ^psi_f[49][7:0];
       end
    100: begin
         out_reg[7:0] <= psi_f[50][15:8];
         parity_reg <= ^psi_f[50][15:8];
       end
    101: begin
         out_reg[7:0] <= psi_f[50][7:0];
         parity_reg <= ^psi_f[50][7:0];
       end
    102: begin
         out_reg[7:0] <= psi_f[51][15:8];
         parity_reg <= ^psi_f[51][15:8];
       end
    103: begin
         out_reg[7:0] <= psi_f[51][7:0];
         parity_reg <= ^psi_f[51][7:0];
       end
    104: begin
         out_reg[7:0] <= psi_f[52][15:8];
         parity_reg <= ^psi_f[52][15:8];
       end
    105: begin
         out_reg[7:0] <= psi_f[52][7:0];
         parity_reg <= ^psi_f[52][7:0];
       end
    106: begin
         out_reg[7:0] <= psi_f[53][15:8];
         parity_reg <= ^psi_f[53][15:8];
       end
    107: begin
         out_reg[7:0] <= psi_f[53][7:0];
         parity_reg <= ^psi_f[53][7:0];
       end
    108: begin
         out_reg[7:0] <= psi_f[54][15:8];
         parity_reg <= ^psi_f[54][15:8];
       end
    109: begin
         out_reg[7:0] <= psi_f[54][7:0];
         parity_reg <= ^psi_f[54][7:0];
       end
    110: begin
         out_reg[7:0] <= psi_f[55][15:8];
         parity_reg <= ^psi_f[55][15:8];
       end
    111: begin
         out_reg[7:0] <= psi_f[55][7:0];
         parity_reg <= ^psi_f[55][7:0];
       end
    112: begin
         out_reg[7:0] <= psi_f[56][15:8];
         parity_reg <= ^psi_f[56][15:8];
       end
    113: begin
         out_reg[7:0] <= psi_f[56][7:0];
         parity_reg <= ^psi_f[56][7:0];
       end
    114: begin
         out_reg[7:0] <= psi_f[57][15:8];
         parity_reg <= ^psi_f[57][15:8];
       end
    115: begin
         out_reg[7:0] <= psi_f[57][7:0];
         parity_reg <= ^psi_f[57][7:0];
       end
    116: begin
         out_reg[7:0] <= psi_f[58][15:8];
         parity_reg <= ^psi_f[58][15:8];
       end
    117: begin
         out_reg[7:0] <= psi_f[58][7:0];
         parity_reg <= ^psi_f[58][7:0];
       end
    118: begin
         out_reg[7:0] <= psi_f[59][15:8];
         parity_reg <= ^psi_f[59][15:8];
       end
    119: begin
         out_reg[7:0] <= psi_f[59][7:0];
         parity_reg <= ^psi_f[59][7:0];
       end
    120: begin
         out_reg[7:0] <= psi_f[60][15:8];
         parity_reg <= ^psi_f[60][15:8];
       end
    121: begin
         out_reg[7:0] <= psi_f[60][7:0];
         parity_reg <= ^psi_f[60][7:0];
       end
    122: begin
         out_reg[7:0] <= psi_f[61][15:8];
         parity_reg <= ^psi_f[61][15:8];
       end
    123: begin
         out_reg[7:0] <= psi_f[61][7:0];
         parity_reg <= ^psi_f[61][7:0];
       end
    124: begin
         out_reg[7:0] <= psi_f[62][15:8];
         parity_reg <= ^psi_f[62][15:8];
       end
    125: begin
         out_reg[7:0] <= psi_f[62][7:0];
         parity_reg <= ^psi_f[62][7:0];
       end
    126: begin
         out_reg[7:0] <= psi_f[63][15:8];
         parity_reg <= ^psi_f[63][15:8];
       end
    127: begin
         out_reg[7:0] <= psi_f[63][7:0];
         parity_reg <= ^psi_f[63][7:0];
       end
    128: begin
         out_reg[7:0] <= psi_f[64][15:8];
         parity_reg <= ^psi_f[64][15:8];
       end
    129: begin
         out_reg[7:0] <= psi_f[64][7:0];
         parity_reg <= ^psi_f[64][7:0];
       end
    130: begin
         out_reg[7:0] <= psi_f[65][15:8];
         parity_reg <= ^psi_f[65][15:8];
       end
    131: begin
         out_reg[7:0] <= psi_f[65][7:0];
         parity_reg <= ^psi_f[65][7:0];
       end
    132: begin
         out_reg[7:0] <= psi_f[66][15:8];
         parity_reg <= ^psi_f[66][15:8];
       end
    133: begin
         out_reg[7:0] <= psi_f[66][7:0];
         parity_reg <= ^psi_f[66][7:0];
       end
    134: begin
         out_reg[7:0] <= psi_f[67][15:8];
         parity_reg <= ^psi_f[67][15:8];
       end
    135: begin
         out_reg[7:0] <= psi_f[67][7:0];
         parity_reg <= ^psi_f[67][7:0];
       end
    136: begin
         out_reg[7:0] <= psi_f[68][15:8];
         parity_reg <= ^psi_f[68][15:8];
       end
    137: begin
         out_reg[7:0] <= psi_f[68][7:0];
         parity_reg <= ^psi_f[68][7:0];
       end
    138: begin
         out_reg[7:0] <= psi_f[69][15:8];
         parity_reg <= ^psi_f[69][15:8];
       end
    139: begin
         out_reg[7:0] <= psi_f[69][7:0];
         parity_reg <= ^psi_f[69][7:0];
       end
    140: begin
         out_reg[7:0] <= psi_f[70][15:8];
         parity_reg <= ^psi_f[70][15:8];
       end
    141: begin
         out_reg[7:0] <= psi_f[70][7:0];
         parity_reg <= ^psi_f[70][7:0];
       end
    142: begin
         out_reg[7:0] <= psi_f[71][15:8];
         parity_reg <= ^psi_f[71][15:8];
       end
    143: begin
         out_reg[7:0] <= psi_f[71][7:0];
         parity_reg <= ^psi_f[71][7:0];
       end
    144: begin
         out_reg[7:0] <= psi_f[72][15:8];
         parity_reg <= ^psi_f[72][15:8];
       end
    145: begin
         out_reg[7:0] <= psi_f[72][7:0];
         parity_reg <= ^psi_f[72][7:0];
       end
    146: begin
         out_reg[7:0] <= psi_f[73][15:8];
         parity_reg <= ^psi_f[73][15:8];
       end
    147: begin
         out_reg[7:0] <= psi_f[73][7:0];
         parity_reg <= ^psi_f[73][7:0];
       end
    148: begin
         out_reg[7:0] <= psi_f[74][15:8];
         parity_reg <= ^psi_f[74][15:8];
       end
    149: begin
         out_reg[7:0] <= psi_f[74][7:0];
         parity_reg <= ^psi_f[74][7:0];
       end
    150: begin
         out_reg[7:0] <= psi_f[75][15:8];
         parity_reg <= ^psi_f[75][15:8];
       end
    151: begin
         out_reg[7:0] <= psi_f[75][7:0];
         parity_reg <= ^psi_f[75][7:0];
       end
    152: begin
         out_reg[7:0] <= psi_f[76][15:8];
         parity_reg <= ^psi_f[76][15:8];
       end
    153: begin
         out_reg[7:0] <= psi_f[76][7:0];
         parity_reg <= ^psi_f[76][7:0];
       end
    154: begin
         out_reg[7:0] <= psi_f[77][15:8];
         parity_reg <= ^psi_f[77][15:8];
       end
    155: begin
         out_reg[7:0] <= psi_f[77][7:0];
         parity_reg <= ^psi_f[77][7:0];
       end
    156: begin
         out_reg[7:0] <= psi_f[78][15:8];
         parity_reg <= ^psi_f[78][15:8];
       end
    157: begin
         out_reg[7:0] <= psi_f[78][7:0];
         parity_reg <= ^psi_f[78][7:0];
       end
    158: begin
         out_reg[7:0] <= psi_f[79][15:8];
         parity_reg <= ^psi_f[79][15:8];
       end
    159: begin
         out_reg[7:0] <= psi_f[79][7:0];
         parity_reg <= ^psi_f[79][7:0];
       end
    160: begin
         out_reg[7:0] <= psi_f[80][15:8];
         parity_reg <= ^psi_f[80][15:8];
       end
    161: begin
         out_reg[7:0] <= psi_f[80][7:0];
         parity_reg <= ^psi_f[80][7:0];
       end
    162: begin
         out_reg[7:0] <= psi_f[81][15:8];
         parity_reg <= ^psi_f[81][15:8];
       end
    163: begin
         out_reg[7:0] <= psi_f[81][7:0];
         parity_reg <= ^psi_f[81][7:0];
       end
    164: begin
         out_reg[7:0] <= psi_f[82][15:8];
         parity_reg <= ^psi_f[82][15:8];
       end
    165: begin
         out_reg[7:0] <= psi_f[82][7:0];
         parity_reg <= ^psi_f[82][7:0];
       end
    166: begin
         out_reg[7:0] <= psi_f[83][15:8];
         parity_reg <= ^psi_f[83][15:8];
       end
    167: begin
         out_reg[7:0] <= psi_f[83][7:0];
         parity_reg <= ^psi_f[83][7:0];
       end
    168: begin
         out_reg[7:0] <= psi_f[84][15:8];
         parity_reg <= ^psi_f[84][15:8];
       end
    169: begin
         out_reg[7:0] <= psi_f[84][7:0];
         parity_reg <= ^psi_f[84][7:0];
       end
    170: begin
         out_reg[7:0] <= psi_f[85][15:8];
         parity_reg <= ^psi_f[85][15:8];
       end
    171: begin
         out_reg[7:0] <= psi_f[85][7:0];
         parity_reg <= ^psi_f[85][7:0];
       end
    172: begin
         out_reg[7:0] <= psi_f[86][15:8];
         parity_reg <= ^psi_f[86][15:8];
       end
    173: begin
         out_reg[7:0] <= psi_f[86][7:0];
         parity_reg <= ^psi_f[86][7:0];
       end
    174: begin
         out_reg[7:0] <= psi_f[87][15:8];
         parity_reg <= ^psi_f[87][15:8];
       end
    175: begin
         out_reg[7:0] <= psi_f[87][7:0];
         parity_reg <= ^psi_f[87][7:0];
       end
    176: begin
         out_reg[7:0] <= psi_f[88][15:8];
         parity_reg <= ^psi_f[88][15:8];
       end
    177: begin
         out_reg[7:0] <= psi_f[88][7:0];
         parity_reg <= ^psi_f[88][7:0];
       end
    178: begin
         out_reg[7:0] <= psi_f[89][15:8];
         parity_reg <= ^psi_f[89][15:8];
       end
    179: begin
         out_reg[7:0] <= psi_f[89][7:0];
         parity_reg <= ^psi_f[89][7:0];
       end
    180: begin
         out_reg[7:0] <= psi_f[90][15:8];
         parity_reg <= ^psi_f[90][15:8];
       end
    181: begin
         out_reg[7:0] <= psi_f[90][7:0];
         parity_reg <= ^psi_f[90][7:0];
       end
    182: begin
         out_reg[7:0] <= psi_f[91][15:8];
         parity_reg <= ^psi_f[91][15:8];
       end
    183: begin
         out_reg[7:0] <= psi_f[91][7:0];
         parity_reg <= ^psi_f[91][7:0];
       end
    184: begin
         out_reg[7:0] <= psi_f[92][15:8];
         parity_reg <= ^psi_f[92][15:8];
       end
    185: begin
         out_reg[7:0] <= psi_f[92][7:0];
         parity_reg <= ^psi_f[92][7:0];
       end
    186: begin
         out_reg[7:0] <= psi_f[93][15:8];
         parity_reg <= ^psi_f[93][15:8];
       end
    187: begin
         out_reg[7:0] <= psi_f[93][7:0];
         parity_reg <= ^psi_f[93][7:0];
       end
    188: begin
         out_reg[7:0] <= psi_f[94][15:8];
         parity_reg <= ^psi_f[94][15:8];
       end
    189: begin
         out_reg[7:0] <= psi_f[94][7:0];
         parity_reg <= ^psi_f[94][7:0];
       end
    190: begin
         out_reg[7:0] <= psi_f[95][15:8];
         parity_reg <= ^psi_f[95][15:8];
       end
    191: begin
         out_reg[7:0] <= psi_f[95][7:0];
         parity_reg <= ^psi_f[95][7:0];
       end
    192: begin
         out_reg[7:0] <= psi_f[96][15:8];
         parity_reg <= ^psi_f[96][15:8];
       end
    193: begin
         out_reg[7:0] <= psi_f[96][7:0];
         parity_reg <= ^psi_f[96][7:0];
       end
    194: begin
         out_reg[7:0] <= psi_f[97][15:8];
         parity_reg <= ^psi_f[97][15:8];
       end
    195: begin
         out_reg[7:0] <= psi_f[97][7:0];
         parity_reg <= ^psi_f[97][7:0];
       end
    196: begin
         out_reg[7:0] <= psi_f[98][15:8];
         parity_reg <= ^psi_f[98][15:8];
       end
    197: begin
         out_reg[7:0] <= psi_f[98][7:0];
         parity_reg <= ^psi_f[98][7:0];
       end
    198: begin
         out_reg[7:0] <= psi_f[99][15:8];
         parity_reg <= ^psi_f[99][15:8];
       end
    199: begin
         out_reg[7:0] <= psi_f[99][7:0];
         parity_reg <= ^psi_f[99][7:0];
       end
    200: begin
         out_reg[7:0] <= psi_f[100][15:8];
         parity_reg <= ^psi_f[100][15:8];
       end
    201: begin
         out_reg[7:0] <= psi_f[100][7:0];
         parity_reg <= ^psi_f[100][7:0];
       end
    202: begin
         out_reg[7:0] <= psi_f[101][15:8];
         parity_reg <= ^psi_f[101][15:8];
       end
    203: begin
         out_reg[7:0] <= psi_f[101][7:0];
         parity_reg <= ^psi_f[101][7:0];
       end
    204: begin
         out_reg[7:0] <= psi_f[102][15:8];
         parity_reg <= ^psi_f[102][15:8];
       end
    205: begin
         out_reg[7:0] <= psi_f[102][7:0];
         parity_reg <= ^psi_f[102][7:0];
       end
    206: begin
         out_reg[7:0] <= psi_f[103][15:8];
         parity_reg <= ^psi_f[103][15:8];
       end
    207: begin
         out_reg[7:0] <= psi_f[103][7:0];
         parity_reg <= ^psi_f[103][7:0];
       end
    208: begin
         out_reg[7:0] <= psi_f[104][15:8];
         parity_reg <= ^psi_f[104][15:8];
       end
    209: begin
         out_reg[7:0] <= psi_f[104][7:0];
         parity_reg <= ^psi_f[104][7:0];
       end
    210: begin
         out_reg[7:0] <= psi_f[105][15:8];
         parity_reg <= ^psi_f[105][15:8];
       end
    211: begin
         out_reg[7:0] <= psi_f[105][7:0];
         parity_reg <= ^psi_f[105][7:0];
       end
    212: begin
         out_reg[7:0] <= psi_f[106][15:8];
         parity_reg <= ^psi_f[106][15:8];
       end
    213: begin
         out_reg[7:0] <= psi_f[106][7:0];
         parity_reg <= ^psi_f[106][7:0];
       end
    214: begin
         out_reg[7:0] <= psi_f[107][15:8];
         parity_reg <= ^psi_f[107][15:8];
       end
    215: begin
         out_reg[7:0] <= psi_f[107][7:0];
         parity_reg <= ^psi_f[107][7:0];
       end
    216: begin
         out_reg[7:0] <= psi_f[108][15:8];
         parity_reg <= ^psi_f[108][15:8];
       end
    217: begin
         out_reg[7:0] <= psi_f[108][7:0];
         parity_reg <= ^psi_f[108][7:0];
       end
    218: begin
         out_reg[7:0] <= psi_f[109][15:8];
         parity_reg <= ^psi_f[109][15:8];
       end
    219: begin
         out_reg[7:0] <= psi_f[109][7:0];
         parity_reg <= ^psi_f[109][7:0];
       end
    220: begin
         out_reg[7:0] <= psi_f[110][15:8];
         parity_reg <= ^psi_f[110][15:8];
       end
    221: begin
         out_reg[7:0] <= psi_f[110][7:0];
         parity_reg <= ^psi_f[110][7:0];
       end
    222: begin
         out_reg[7:0] <= psi_f[111][15:8];
         parity_reg <= ^psi_f[111][15:8];
       end
    223: begin
         out_reg[7:0] <= psi_f[111][7:0];
         parity_reg <= ^psi_f[111][7:0];
       end
    224: begin
         out_reg[7:0] <= psi_f[112][15:8];
         parity_reg <= ^psi_f[112][15:8];
       end
    225: begin
         out_reg[7:0] <= psi_f[112][7:0];
         parity_reg <= ^psi_f[112][7:0];
       end
    226: begin
         out_reg[7:0] <= psi_f[113][15:8];
         parity_reg <= ^psi_f[113][15:8];
       end
    227: begin
         out_reg[7:0] <= psi_f[113][7:0];
         parity_reg <= ^psi_f[113][7:0];
       end
    228: begin
         out_reg[7:0] <= psi_f[114][15:8];
         parity_reg <= ^psi_f[114][15:8];
       end
    229: begin
         out_reg[7:0] <= psi_f[114][7:0];
         parity_reg <= ^psi_f[114][7:0];
       end
    230: begin
         out_reg[7:0] <= psi_f[115][15:8];
         parity_reg <= ^psi_f[115][15:8];
       end
    231: begin
         out_reg[7:0] <= psi_f[115][7:0];
         parity_reg <= ^psi_f[115][7:0];
       end
    232: begin
         out_reg[7:0] <= psi_f[116][15:8];
         parity_reg <= ^psi_f[116][15:8];
       end
    233: begin
         out_reg[7:0] <= psi_f[116][7:0];
         parity_reg <= ^psi_f[116][7:0];
       end
    234: begin
         out_reg[7:0] <= psi_f[117][15:8];
         parity_reg <= ^psi_f[117][15:8];
       end
    235: begin
         out_reg[7:0] <= psi_f[117][7:0];
         parity_reg <= ^psi_f[117][7:0];
       end
    236: begin
         out_reg[7:0] <= psi_f[118][15:8];
         parity_reg <= ^psi_f[118][15:8];
       end
    237: begin
         out_reg[7:0] <= psi_f[118][7:0];
         parity_reg <= ^psi_f[118][7:0];
       end
    238: begin
         out_reg[7:0] <= psi_f[119][15:8];
         parity_reg <= ^psi_f[119][15:8];
       end
    239: begin
         out_reg[7:0] <= psi_f[119][7:0];
         parity_reg <= ^psi_f[119][7:0];
       end
    240: begin
         out_reg[7:0] <= psi_f[120][15:8];
         parity_reg <= ^psi_f[120][15:8];
       end
    241: begin
         out_reg[7:0] <= psi_f[120][7:0];
         parity_reg <= ^psi_f[120][7:0];
       end
    242: begin
         out_reg[7:0] <= psi_f[121][15:8];
         parity_reg <= ^psi_f[121][15:8];
       end
    243: begin
         out_reg[7:0] <= psi_f[121][7:0];
         parity_reg <= ^psi_f[121][7:0];
       end
    244: begin
         out_reg[7:0] <= psi_f[122][15:8];
         parity_reg <= ^psi_f[122][15:8];
       end
    245: begin
         out_reg[7:0] <= psi_f[122][7:0];
         parity_reg <= ^psi_f[122][7:0];
       end
    246: begin
         out_reg[7:0] <= psi_f[123][15:8];
         parity_reg <= ^psi_f[123][15:8];
       end
    247: begin
         out_reg[7:0] <= psi_f[123][7:0];
         parity_reg <= ^psi_f[123][7:0];
       end
    248: begin
         out_reg[7:0] <= psi_f[124][15:8];
         parity_reg <= ^psi_f[124][15:8];
       end
    249: begin
         out_reg[7:0] <= psi_f[124][7:0];
         parity_reg <= ^psi_f[124][7:0];
       end
    250: begin
         out_reg[7:0] <= psi_f[125][15:8];
         parity_reg <= ^psi_f[125][15:8];
       end
    251: begin
         out_reg[7:0] <= psi_f[125][7:0];
         parity_reg <= ^psi_f[125][7:0];
       end
    252: begin
         out_reg[7:0] <= psi_f[126][15:8];
         parity_reg <= ^psi_f[126][15:8];
       end
    253: begin
         out_reg[7:0] <= psi_f[126][7:0];
         parity_reg <= ^psi_f[126][7:0];
       end
    254: begin
         out_reg[7:0] <= psi_f[127][15:8];
         parity_reg <= ^psi_f[127][15:8];
       end
    255: begin
         out_reg[7:0] <= psi_f[127][7:0];
         parity_reg <= ^psi_f[127][7:0];
       end
    256: begin
         out_reg[7:0] <= psi_f[128][15:8];
         parity_reg <= ^psi_f[128][15:8];
       end
    257: begin
         out_reg[7:0] <= psi_f[128][7:0];
         parity_reg <= ^psi_f[128][7:0];
       end
    258: begin
         out_reg[7:0] <= psi_f[129][15:8];
         parity_reg <= ^psi_f[129][15:8];
       end
    259: begin
         out_reg[7:0] <= psi_f[129][7:0];
         parity_reg <= ^psi_f[129][7:0];
       end
    260: begin
         out_reg[7:0] <= psi_f[130][15:8];
         parity_reg <= ^psi_f[130][15:8];
       end
    261: begin
         out_reg[7:0] <= psi_f[130][7:0];
         parity_reg <= ^psi_f[130][7:0];
       end
    262: begin
         out_reg[7:0] <= psi_f[131][15:8];
         parity_reg <= ^psi_f[131][15:8];
       end
    263: begin
         out_reg[7:0] <= psi_f[131][7:0];
         parity_reg <= ^psi_f[131][7:0];
       end
    264: begin
         out_reg[7:0] <= psi_f[132][15:8];
         parity_reg <= ^psi_f[132][15:8];
       end
    265: begin
         out_reg[7:0] <= psi_f[132][7:0];
         parity_reg <= ^psi_f[132][7:0];
       end
    266: begin
         out_reg[7:0] <= psi_f[133][15:8];
         parity_reg <= ^psi_f[133][15:8];
       end
    267: begin
         out_reg[7:0] <= psi_f[133][7:0];
         parity_reg <= ^psi_f[133][7:0];
       end
    268: begin
         out_reg[7:0] <= psi_f[134][15:8];
         parity_reg <= ^psi_f[134][15:8];
       end
    269: begin
         out_reg[7:0] <= psi_f[134][7:0];
         parity_reg <= ^psi_f[134][7:0];
       end
    270: begin
         out_reg[7:0] <= psi_f[135][15:8];
         parity_reg <= ^psi_f[135][15:8];
       end
    271: begin
         out_reg[7:0] <= psi_f[135][7:0];
         parity_reg <= ^psi_f[135][7:0];
       end
    272: begin
         out_reg[7:0] <= psi_f[136][15:8];
         parity_reg <= ^psi_f[136][15:8];
       end
    273: begin
         out_reg[7:0] <= psi_f[136][7:0];
         parity_reg <= ^psi_f[136][7:0];
       end
    274: begin
         out_reg[7:0] <= psi_f[137][15:8];
         parity_reg <= ^psi_f[137][15:8];
       end
    275: begin
         out_reg[7:0] <= psi_f[137][7:0];
         parity_reg <= ^psi_f[137][7:0];
       end
    276: begin
         out_reg[7:0] <= psi_f[138][15:8];
         parity_reg <= ^psi_f[138][15:8];
       end
    277: begin
         out_reg[7:0] <= psi_f[138][7:0];
         parity_reg <= ^psi_f[138][7:0];
       end
    278: begin
         out_reg[7:0] <= psi_f[139][15:8];
         parity_reg <= ^psi_f[139][15:8];
       end
    279: begin
         out_reg[7:0] <= psi_f[139][7:0];
         parity_reg <= ^psi_f[139][7:0];
       end
    280: begin
         out_reg[7:0] <= psi_f[140][15:8];
         parity_reg <= ^psi_f[140][15:8];
       end
    281: begin
         out_reg[7:0] <= psi_f[140][7:0];
         parity_reg <= ^psi_f[140][7:0];
       end
    282: begin
         out_reg[7:0] <= psi_f[141][15:8];
         parity_reg <= ^psi_f[141][15:8];
       end
    283: begin
         out_reg[7:0] <= psi_f[141][7:0];
         parity_reg <= ^psi_f[141][7:0];
       end
    284: begin
         out_reg[7:0] <= psi_f[142][15:8];
         parity_reg <= ^psi_f[142][15:8];
       end
    285: begin
         out_reg[7:0] <= psi_f[142][7:0];
         parity_reg <= ^psi_f[142][7:0];
       end
    286: begin
         out_reg[7:0] <= psi_f[143][15:8];
         parity_reg <= ^psi_f[143][15:8];
       end
    287: begin
         out_reg[7:0] <= psi_f[143][7:0];
         parity_reg <= ^psi_f[143][7:0];
       end
    288: begin
         out_reg[7:0] <= psi_f[144][15:8];
         parity_reg <= ^psi_f[144][15:8];
       end
    289: begin
         out_reg[7:0] <= psi_f[144][7:0];
         parity_reg <= ^psi_f[144][7:0];
       end
    290: begin
         out_reg[7:0] <= psi_f[145][15:8];
         parity_reg <= ^psi_f[145][15:8];
       end
    291: begin
         out_reg[7:0] <= psi_f[145][7:0];
         parity_reg <= ^psi_f[145][7:0];
       end
    292: begin
         out_reg[7:0] <= psi_f[146][15:8];
         parity_reg <= ^psi_f[146][15:8];
       end
    293: begin
         out_reg[7:0] <= psi_f[146][7:0];
         parity_reg <= ^psi_f[146][7:0];
       end
    294: begin
         out_reg[7:0] <= psi_f[147][15:8];
         parity_reg <= ^psi_f[147][15:8];
       end
    295: begin
         out_reg[7:0] <= psi_f[147][7:0];
         parity_reg <= ^psi_f[147][7:0];
       end
    296: begin
         out_reg[7:0] <= psi_f[148][15:8];
         parity_reg <= ^psi_f[148][15:8];
       end
    297: begin
         out_reg[7:0] <= psi_f[148][7:0];
         parity_reg <= ^psi_f[148][7:0];
       end
    298: begin
         out_reg[7:0] <= psi_f[149][15:8];
         parity_reg <= ^psi_f[149][15:8];
       end
    299: begin
         out_reg[7:0] <= psi_f[149][7:0];
         parity_reg <= ^psi_f[149][7:0];
       end
    300: begin
         out_reg[7:0] <= psi_f[150][15:8];
         parity_reg <= ^psi_f[150][15:8];
       end
    301: begin
         out_reg[7:0] <= psi_f[150][7:0];
         parity_reg <= ^psi_f[150][7:0];
       end
    302: begin
         out_reg[7:0] <= psi_f[151][15:8];
         parity_reg <= ^psi_f[151][15:8];
       end
    303: begin
         out_reg[7:0] <= psi_f[151][7:0];
         parity_reg <= ^psi_f[151][7:0];
       end
    304: begin
         out_reg[7:0] <= psi_f[152][15:8];
         parity_reg <= ^psi_f[152][15:8];
       end
    305: begin
         out_reg[7:0] <= psi_f[152][7:0];
         parity_reg <= ^psi_f[152][7:0];
       end
    306: begin
         out_reg[7:0] <= psi_f[153][15:8];
         parity_reg <= ^psi_f[153][15:8];
       end
    307: begin
         out_reg[7:0] <= psi_f[153][7:0];
         parity_reg <= ^psi_f[153][7:0];
       end
    308: begin
         out_reg[7:0] <= psi_f[154][15:8];
         parity_reg <= ^psi_f[154][15:8];
       end
    309: begin
         out_reg[7:0] <= psi_f[154][7:0];
         parity_reg <= ^psi_f[154][7:0];
       end
    310: begin
         out_reg[7:0] <= psi_f[155][15:8];
         parity_reg <= ^psi_f[155][15:8];
       end
    311: begin
         out_reg[7:0] <= psi_f[155][7:0];
         parity_reg <= ^psi_f[155][7:0];
       end
    312: begin
         out_reg[7:0] <= psi_f[156][15:8];
         parity_reg <= ^psi_f[156][15:8];
       end
    313: begin
         out_reg[7:0] <= psi_f[156][7:0];
         parity_reg <= ^psi_f[156][7:0];
       end
    314: begin
         out_reg[7:0] <= psi_f[157][15:8];
         parity_reg <= ^psi_f[157][15:8];
       end
    315: begin
         out_reg[7:0] <= psi_f[157][7:0];
         parity_reg <= ^psi_f[157][7:0];
       end
    316: begin
         out_reg[7:0] <= psi_f[158][15:8];
         parity_reg <= ^psi_f[158][15:8];
       end
    317: begin
         out_reg[7:0] <= psi_f[158][7:0];
         parity_reg <= ^psi_f[158][7:0];
       end
    318: begin
         out_reg[7:0] <= psi_f[159][15:8];
         parity_reg <= ^psi_f[159][15:8];
       end
    319: begin
         out_reg[7:0] <= psi_f[159][7:0];
         parity_reg <= ^psi_f[159][7:0];
       end
    320: begin
         out_reg[7:0] <= psi_f[160][15:8];
         parity_reg <= ^psi_f[160][15:8];
       end
    321: begin
         out_reg[7:0] <= psi_f[160][7:0];
         parity_reg <= ^psi_f[160][7:0];
       end
    322: begin
         out_reg[7:0] <= psi_f[161][15:8];
         parity_reg <= ^psi_f[161][15:8];
       end
    323: begin
         out_reg[7:0] <= psi_f[161][7:0];
         parity_reg <= ^psi_f[161][7:0];
       end
    324: begin
         out_reg[7:0] <= psi_f[162][15:8];
         parity_reg <= ^psi_f[162][15:8];
       end
    325: begin
         out_reg[7:0] <= psi_f[162][7:0];
         parity_reg <= ^psi_f[162][7:0];
       end
    326: begin
         out_reg[7:0] <= psi_f[163][15:8];
         parity_reg <= ^psi_f[163][15:8];
       end
    327: begin
         out_reg[7:0] <= psi_f[163][7:0];
         parity_reg <= ^psi_f[163][7:0];
       end
    328: begin
         out_reg[7:0] <= psi_f[164][15:8];
         parity_reg <= ^psi_f[164][15:8];
       end
    329: begin
         out_reg[7:0] <= psi_f[164][7:0];
         parity_reg <= ^psi_f[164][7:0];
       end
    330: begin
         out_reg[7:0] <= psi_f[165][15:8];
         parity_reg <= ^psi_f[165][15:8];
       end
    331: begin
         out_reg[7:0] <= psi_f[165][7:0];
         parity_reg <= ^psi_f[165][7:0];
       end
    332: begin
         out_reg[7:0] <= psi_f[166][15:8];
         parity_reg <= ^psi_f[166][15:8];
       end
    333: begin
         out_reg[7:0] <= psi_f[166][7:0];
         parity_reg <= ^psi_f[166][7:0];
       end
    334: begin
         out_reg[7:0] <= psi_f[167][15:8];
         parity_reg <= ^psi_f[167][15:8];
       end
    335: begin
         out_reg[7:0] <= psi_f[167][7:0];
         parity_reg <= ^psi_f[167][7:0];
       end
    336: begin
         out_reg[7:0] <= psi_f[168][15:8];
         parity_reg <= ^psi_f[168][15:8];
       end
    337: begin
         out_reg[7:0] <= psi_f[168][7:0];
         parity_reg <= ^psi_f[168][7:0];
       end
    338: begin
         out_reg[7:0] <= psi_f[169][15:8];
         parity_reg <= ^psi_f[169][15:8];
       end
    339: begin
         out_reg[7:0] <= psi_f[169][7:0];
         parity_reg <= ^psi_f[169][7:0];
       end
    340: begin
         out_reg[7:0] <= psi_f[170][15:8];
         parity_reg <= ^psi_f[170][15:8];
       end
    341: begin
         out_reg[7:0] <= psi_f[170][7:0];
         parity_reg <= ^psi_f[170][7:0];
       end
    342: begin
         out_reg[7:0] <= psi_f[171][15:8];
         parity_reg <= ^psi_f[171][15:8];
       end
    343: begin
         out_reg[7:0] <= psi_f[171][7:0];
         parity_reg <= ^psi_f[171][7:0];
       end
    344: begin
         out_reg[7:0] <= psi_f[172][15:8];
         parity_reg <= ^psi_f[172][15:8];
       end
    345: begin
         out_reg[7:0] <= psi_f[172][7:0];
         parity_reg <= ^psi_f[172][7:0];
       end
    346: begin
         out_reg[7:0] <= psi_f[173][15:8];
         parity_reg <= ^psi_f[173][15:8];
       end
    347: begin
         out_reg[7:0] <= psi_f[173][7:0];
         parity_reg <= ^psi_f[173][7:0];
       end
    348: begin
         out_reg[7:0] <= psi_f[174][15:8];
         parity_reg <= ^psi_f[174][15:8];
       end
    349: begin
         out_reg[7:0] <= psi_f[174][7:0];
         parity_reg <= ^psi_f[174][7:0];
       end
    350: begin
         out_reg[7:0] <= psi_f[175][15:8];
         parity_reg <= ^psi_f[175][15:8];
       end
    351: begin
         out_reg[7:0] <= psi_f[175][7:0];
         parity_reg <= ^psi_f[175][7:0];
       end
    352: begin
         out_reg[7:0] <= psi_f[176][15:8];
         parity_reg <= ^psi_f[176][15:8];
       end
    353: begin
         out_reg[7:0] <= psi_f[176][7:0];
         parity_reg <= ^psi_f[176][7:0];
       end
    354: begin
         out_reg[7:0] <= psi_f[177][15:8];
         parity_reg <= ^psi_f[177][15:8];
       end
    355: begin
         out_reg[7:0] <= psi_f[177][7:0];
         parity_reg <= ^psi_f[177][7:0];
       end
    356: begin
         out_reg[7:0] <= psi_f[178][15:8];
         parity_reg <= ^psi_f[178][15:8];
       end
    357: begin
         out_reg[7:0] <= psi_f[178][7:0];
         parity_reg <= ^psi_f[178][7:0];
       end
    358: begin
         out_reg[7:0] <= psi_f[179][15:8];
         parity_reg <= ^psi_f[179][15:8];
       end
    359: begin
         out_reg[7:0] <= psi_f[179][7:0];
         parity_reg <= ^psi_f[179][7:0];
       end
    360: begin
         out_reg[7:0] <= psi_f[180][15:8];
         parity_reg <= ^psi_f[180][15:8];
       end
    361: begin
         out_reg[7:0] <= psi_f[180][7:0];
         parity_reg <= ^psi_f[180][7:0];
       end
    362: begin
         out_reg[7:0] <= psi_f[181][15:8];
         parity_reg <= ^psi_f[181][15:8];
       end
    363: begin
         out_reg[7:0] <= psi_f[181][7:0];
         parity_reg <= ^psi_f[181][7:0];
       end
    364: begin
         out_reg[7:0] <= psi_f[182][15:8];
         parity_reg <= ^psi_f[182][15:8];
       end
    365: begin
         out_reg[7:0] <= psi_f[182][7:0];
         parity_reg <= ^psi_f[182][7:0];
       end
    366: begin
         out_reg[7:0] <= psi_f[183][15:8];
         parity_reg <= ^psi_f[183][15:8];
       end
    367: begin
         out_reg[7:0] <= psi_f[183][7:0];
         parity_reg <= ^psi_f[183][7:0];
       end
    368: begin
         out_reg[7:0] <= psi_f[184][15:8];
         parity_reg <= ^psi_f[184][15:8];
       end
    369: begin
         out_reg[7:0] <= psi_f[184][7:0];
         parity_reg <= ^psi_f[184][7:0];
       end
    370: begin
         out_reg[7:0] <= psi_f[185][15:8];
         parity_reg <= ^psi_f[185][15:8];
       end
    371: begin
         out_reg[7:0] <= psi_f[185][7:0];
         parity_reg <= ^psi_f[185][7:0];
       end
    372: begin
         out_reg[7:0] <= psi_f[186][15:8];
         parity_reg <= ^psi_f[186][15:8];
       end
    373: begin
         out_reg[7:0] <= psi_f[186][7:0];
         parity_reg <= ^psi_f[186][7:0];
       end
    374: begin
         out_reg[7:0] <= psi_f[187][15:8];
         parity_reg <= ^psi_f[187][15:8];
       end
    375: begin
         out_reg[7:0] <= psi_f[187][7:0];
         parity_reg <= ^psi_f[187][7:0];
       end
    376: begin
         out_reg[7:0] <= psi_f[188][15:8];
         parity_reg <= ^psi_f[188][15:8];
       end
    377: begin
         out_reg[7:0] <= psi_f[188][7:0];
         parity_reg <= ^psi_f[188][7:0];
       end
    378: begin
         out_reg[7:0] <= psi_f[189][15:8];
         parity_reg <= ^psi_f[189][15:8];
       end
    379: begin
         out_reg[7:0] <= psi_f[189][7:0];
         parity_reg <= ^psi_f[189][7:0];
       end
    380: begin
         out_reg[7:0] <= psi_f[190][15:8];
         parity_reg <= ^psi_f[190][15:8];
       end
    381: begin
         out_reg[7:0] <= psi_f[190][7:0];
         parity_reg <= ^psi_f[190][7:0];
       end
    382: begin
         out_reg[7:0] <= psi_f[191][15:8];
         parity_reg <= ^psi_f[191][15:8];
       end
    383: begin
         out_reg[7:0] <= psi_f[191][7:0];
         parity_reg <= ^psi_f[191][7:0];
       end
    384: begin
         out_reg[7:0] <= psi_f[192][15:8];
         parity_reg <= ^psi_f[192][15:8];
       end
    385: begin
         out_reg[7:0] <= psi_f[192][7:0];
         parity_reg <= ^psi_f[192][7:0];
       end
    386: begin
         out_reg[7:0] <= psi_f[193][15:8];
         parity_reg <= ^psi_f[193][15:8];
       end
    387: begin
         out_reg[7:0] <= psi_f[193][7:0];
         parity_reg <= ^psi_f[193][7:0];
       end
    388: begin
         out_reg[7:0] <= psi_f[194][15:8];
         parity_reg <= ^psi_f[194][15:8];
       end
    389: begin
         out_reg[7:0] <= psi_f[194][7:0];
         parity_reg <= ^psi_f[194][7:0];
       end
    390: begin
         out_reg[7:0] <= psi_f[195][15:8];
         parity_reg <= ^psi_f[195][15:8];
       end
    391: begin
         out_reg[7:0] <= psi_f[195][7:0];
         parity_reg <= ^psi_f[195][7:0];
       end
    392: begin
         out_reg[7:0] <= psi_f[196][15:8];
         parity_reg <= ^psi_f[196][15:8];
       end
    393: begin
         out_reg[7:0] <= psi_f[196][7:0];
         parity_reg <= ^psi_f[196][7:0];
       end
    394: begin
         out_reg[7:0] <= psi_f[197][15:8];
         parity_reg <= ^psi_f[197][15:8];
       end
    395: begin
         out_reg[7:0] <= psi_f[197][7:0];
         parity_reg <= ^psi_f[197][7:0];
       end
    396: begin
         out_reg[7:0] <= psi_f[198][15:8];
         parity_reg <= ^psi_f[198][15:8];
       end
    397: begin
         out_reg[7:0] <= psi_f[198][7:0];
         parity_reg <= ^psi_f[198][7:0];
       end
    398: begin
         out_reg[7:0] <= psi_f[199][15:8];
         parity_reg <= ^psi_f[199][15:8];
       end
    399: begin
         out_reg[7:0] <= psi_f[199][7:0];
         parity_reg <= ^psi_f[199][7:0];
       end
    400: begin
         out_reg[7:0] <= psi_f[200][15:8];
         parity_reg <= ^psi_f[200][15:8];
       end
    401: begin
         out_reg[7:0] <= psi_f[200][7:0];
         parity_reg <= ^psi_f[200][7:0];
       end
    402: begin
         out_reg[7:0] <= psi_f[201][15:8];
         parity_reg <= ^psi_f[201][15:8];
       end
    403: begin
         out_reg[7:0] <= psi_f[201][7:0];
         parity_reg <= ^psi_f[201][7:0];
       end
    404: begin
         out_reg[7:0] <= psi_f[202][15:8];
         parity_reg <= ^psi_f[202][15:8];
       end
    405: begin
         out_reg[7:0] <= psi_f[202][7:0];
         parity_reg <= ^psi_f[202][7:0];
       end
    406: begin
         out_reg[7:0] <= psi_f[203][15:8];
         parity_reg <= ^psi_f[203][15:8];
       end
    407: begin
         out_reg[7:0] <= psi_f[203][7:0];
         parity_reg <= ^psi_f[203][7:0];
       end
    408: begin
         out_reg[7:0] <= psi_f[204][15:8];
         parity_reg <= ^psi_f[204][15:8];
       end
    409: begin
         out_reg[7:0] <= psi_f[204][7:0];
         parity_reg <= ^psi_f[204][7:0];
       end
    410: begin
         out_reg[7:0] <= psi_f[205][15:8];
         parity_reg <= ^psi_f[205][15:8];
       end
    411: begin
         out_reg[7:0] <= psi_f[205][7:0];
         parity_reg <= ^psi_f[205][7:0];
       end
    412: begin
         out_reg[7:0] <= psi_f[206][15:8];
         parity_reg <= ^psi_f[206][15:8];
       end
    413: begin
         out_reg[7:0] <= psi_f[206][7:0];
         parity_reg <= ^psi_f[206][7:0];
       end
    414: begin
         out_reg[7:0] <= psi_f[207][15:8];
         parity_reg <= ^psi_f[207][15:8];
       end
    415: begin
         out_reg[7:0] <= psi_f[207][7:0];
         parity_reg <= ^psi_f[207][7:0];
       end
    416: begin
         out_reg[7:0] <= psi_f[208][15:8];
         parity_reg <= ^psi_f[208][15:8];
       end
    417: begin
         out_reg[7:0] <= psi_f[208][7:0];
         parity_reg <= ^psi_f[208][7:0];
       end
    418: begin
         out_reg[7:0] <= psi_f[209][15:8];
         parity_reg <= ^psi_f[209][15:8];
       end
    419: begin
         out_reg[7:0] <= psi_f[209][7:0];
         parity_reg <= ^psi_f[209][7:0];
       end
    420: begin
         out_reg[7:0] <= psi_f[210][15:8];
         parity_reg <= ^psi_f[210][15:8];
       end
    421: begin
         out_reg[7:0] <= psi_f[210][7:0];
         parity_reg <= ^psi_f[210][7:0];
       end
    422: begin
         out_reg[7:0] <= psi_f[211][15:8];
         parity_reg <= ^psi_f[211][15:8];
       end
    423: begin
         out_reg[7:0] <= psi_f[211][7:0];
         parity_reg <= ^psi_f[211][7:0];
       end
    424: begin
         out_reg[7:0] <= psi_f[212][15:8];
         parity_reg <= ^psi_f[212][15:8];
       end
    425: begin
         out_reg[7:0] <= psi_f[212][7:0];
         parity_reg <= ^psi_f[212][7:0];
       end
    426: begin
         out_reg[7:0] <= psi_f[213][15:8];
         parity_reg <= ^psi_f[213][15:8];
       end
    427: begin
         out_reg[7:0] <= psi_f[213][7:0];
         parity_reg <= ^psi_f[213][7:0];
       end
    428: begin
         out_reg[7:0] <= psi_f[214][15:8];
         parity_reg <= ^psi_f[214][15:8];
       end
    429: begin
         out_reg[7:0] <= psi_f[214][7:0];
         parity_reg <= ^psi_f[214][7:0];
       end
    430: begin
         out_reg[7:0] <= psi_f[215][15:8];
         parity_reg <= ^psi_f[215][15:8];
       end
    431: begin
         out_reg[7:0] <= psi_f[215][7:0];
         parity_reg <= ^psi_f[215][7:0];
       end
    432: begin
         out_reg[7:0] <= psi_f[216][15:8];
         parity_reg <= ^psi_f[216][15:8];
       end
    433: begin
         out_reg[7:0] <= psi_f[216][7:0];
         parity_reg <= ^psi_f[216][7:0];
       end
    434: begin
         out_reg[7:0] <= psi_f[217][15:8];
         parity_reg <= ^psi_f[217][15:8];
       end
    435: begin
         out_reg[7:0] <= psi_f[217][7:0];
         parity_reg <= ^psi_f[217][7:0];
       end
    436: begin
         out_reg[7:0] <= psi_f[218][15:8];
         parity_reg <= ^psi_f[218][15:8];
       end
    437: begin
         out_reg[7:0] <= psi_f[218][7:0];
         parity_reg <= ^psi_f[218][7:0];
       end
    438: begin
         out_reg[7:0] <= psi_f[219][15:8];
         parity_reg <= ^psi_f[219][15:8];
       end
    439: begin
         out_reg[7:0] <= psi_f[219][7:0];
         parity_reg <= ^psi_f[219][7:0];
       end
    440: begin
         out_reg[7:0] <= psi_f[220][15:8];
         parity_reg <= ^psi_f[220][15:8];
       end
    441: begin
         out_reg[7:0] <= psi_f[220][7:0];
         parity_reg <= ^psi_f[220][7:0];
       end
    442: begin
         out_reg[7:0] <= psi_f[221][15:8];
         parity_reg <= ^psi_f[221][15:8];
       end
    443: begin
         out_reg[7:0] <= psi_f[221][7:0];
         parity_reg <= ^psi_f[221][7:0];
       end
    444: begin
         out_reg[7:0] <= psi_f[222][15:8];
         parity_reg <= ^psi_f[222][15:8];
       end
    445: begin
         out_reg[7:0] <= psi_f[222][7:0];
         parity_reg <= ^psi_f[222][7:0];
       end
    446: begin
         out_reg[7:0] <= psi_f[223][15:8];
         parity_reg <= ^psi_f[223][15:8];
       end
    447: begin
         out_reg[7:0] <= psi_f[223][7:0];
         parity_reg <= ^psi_f[223][7:0];
       end
    448: begin
         out_reg[7:0] <= psi_f[224][15:8];
         parity_reg <= ^psi_f[224][15:8];
       end
    449: begin
         out_reg[7:0] <= psi_f[224][7:0];
         parity_reg <= ^psi_f[224][7:0];
       end
    450: begin
         out_reg[7:0] <= psi_f[225][15:8];
         parity_reg <= ^psi_f[225][15:8];
       end
    451: begin
         out_reg[7:0] <= psi_f[225][7:0];
         parity_reg <= ^psi_f[225][7:0];
       end
    452: begin
         out_reg[7:0] <= psi_f[226][15:8];
         parity_reg <= ^psi_f[226][15:8];
       end
    453: begin
         out_reg[7:0] <= psi_f[226][7:0];
         parity_reg <= ^psi_f[226][7:0];
       end
    454: begin
         out_reg[7:0] <= psi_f[227][15:8];
         parity_reg <= ^psi_f[227][15:8];
       end
    455: begin
         out_reg[7:0] <= psi_f[227][7:0];
         parity_reg <= ^psi_f[227][7:0];
       end
    456: begin
         out_reg[7:0] <= psi_f[228][15:8];
         parity_reg <= ^psi_f[228][15:8];
       end
    457: begin
         out_reg[7:0] <= psi_f[228][7:0];
         parity_reg <= ^psi_f[228][7:0];
       end
    458: begin
         out_reg[7:0] <= psi_f[229][15:8];
         parity_reg <= ^psi_f[229][15:8];
       end
    459: begin
         out_reg[7:0] <= psi_f[229][7:0];
         parity_reg <= ^psi_f[229][7:0];
       end
    460: begin
         out_reg[7:0] <= psi_f[230][15:8];
         parity_reg <= ^psi_f[230][15:8];
       end
    461: begin
         out_reg[7:0] <= psi_f[230][7:0];
         parity_reg <= ^psi_f[230][7:0];
       end
    462: begin
         out_reg[7:0] <= psi_f[231][15:8];
         parity_reg <= ^psi_f[231][15:8];
       end
    463: begin
         out_reg[7:0] <= psi_f[231][7:0];
         parity_reg <= ^psi_f[231][7:0];
       end
    464: begin
         out_reg[7:0] <= psi_f[232][15:8];
         parity_reg <= ^psi_f[232][15:8];
       end
    465: begin
         out_reg[7:0] <= psi_f[232][7:0];
         parity_reg <= ^psi_f[232][7:0];
       end
    466: begin
         out_reg[7:0] <= psi_f[233][15:8];
         parity_reg <= ^psi_f[233][15:8];
       end
    467: begin
         out_reg[7:0] <= psi_f[233][7:0];
         parity_reg <= ^psi_f[233][7:0];
       end
    468: begin
         out_reg[7:0] <= psi_f[234][15:8];
         parity_reg <= ^psi_f[234][15:8];
       end
    469: begin
         out_reg[7:0] <= psi_f[234][7:0];
         parity_reg <= ^psi_f[234][7:0];
       end
    470: begin
         out_reg[7:0] <= psi_f[235][15:8];
         parity_reg <= ^psi_f[235][15:8];
       end
    471: begin
         out_reg[7:0] <= psi_f[235][7:0];
         parity_reg <= ^psi_f[235][7:0];
       end
    472: begin
         out_reg[7:0] <= psi_f[236][15:8];
         parity_reg <= ^psi_f[236][15:8];
       end
    473: begin
         out_reg[7:0] <= psi_f[236][7:0];
         parity_reg <= ^psi_f[236][7:0];
       end
    474: begin
         out_reg[7:0] <= psi_f[237][15:8];
         parity_reg <= ^psi_f[237][15:8];
       end
    475: begin
         out_reg[7:0] <= psi_f[237][7:0];
         parity_reg <= ^psi_f[237][7:0];
       end
    476: begin
         out_reg[7:0] <= psi_f[238][15:8];
         parity_reg <= ^psi_f[238][15:8];
       end
    477: begin
         out_reg[7:0] <= psi_f[238][7:0];
         parity_reg <= ^psi_f[238][7:0];
       end
    478: begin
         out_reg[7:0] <= psi_f[239][15:8];
         parity_reg <= ^psi_f[239][15:8];
       end
    479: begin
         out_reg[7:0] <= psi_f[239][7:0];
         parity_reg <= ^psi_f[239][7:0];
       end
    480: begin
         out_reg[7:0] <= psi_f[240][15:8];
         parity_reg <= ^psi_f[240][15:8];
       end
    481: begin
         out_reg[7:0] <= psi_f[240][7:0];
         parity_reg <= ^psi_f[240][7:0];
       end
    482: begin
         out_reg[7:0] <= psi_f[241][15:8];
         parity_reg <= ^psi_f[241][15:8];
       end
    483: begin
         out_reg[7:0] <= psi_f[241][7:0];
         parity_reg <= ^psi_f[241][7:0];
       end
    484: begin
         out_reg[7:0] <= psi_f[242][15:8];
         parity_reg <= ^psi_f[242][15:8];
       end
    485: begin
         out_reg[7:0] <= psi_f[242][7:0];
         parity_reg <= ^psi_f[242][7:0];
       end
    486: begin
         out_reg[7:0] <= psi_f[243][15:8];
         parity_reg <= ^psi_f[243][15:8];
       end
    487: begin
         out_reg[7:0] <= psi_f[243][7:0];
         parity_reg <= ^psi_f[243][7:0];
       end
    488: begin
         out_reg[7:0] <= psi_f[244][15:8];
         parity_reg <= ^psi_f[244][15:8];
       end
    489: begin
         out_reg[7:0] <= psi_f[244][7:0];
         parity_reg <= ^psi_f[244][7:0];
       end
    490: begin
         out_reg[7:0] <= psi_f[245][15:8];
         parity_reg <= ^psi_f[245][15:8];
       end
    491: begin
         out_reg[7:0] <= psi_f[245][7:0];
         parity_reg <= ^psi_f[245][7:0];
       end
    492: begin
         out_reg[7:0] <= psi_f[246][15:8];
         parity_reg <= ^psi_f[246][15:8];
       end
    493: begin
         out_reg[7:0] <= psi_f[246][7:0];
         parity_reg <= ^psi_f[246][7:0];
       end
    494: begin
         out_reg[7:0] <= psi_f[247][15:8];
         parity_reg <= ^psi_f[247][15:8];
       end
    495: begin
         out_reg[7:0] <= psi_f[247][7:0];
         parity_reg <= ^psi_f[247][7:0];
       end
    496: begin
         out_reg[7:0] <= psi_f[248][15:8];
         parity_reg <= ^psi_f[248][15:8];
       end
    497: begin
         out_reg[7:0] <= psi_f[248][7:0];
         parity_reg <= ^psi_f[248][7:0];
       end
    498: begin
         out_reg[7:0] <= psi_f[249][15:8];
         parity_reg <= ^psi_f[249][15:8];
       end
    499: begin
         out_reg[7:0] <= psi_f[249][7:0];
         parity_reg <= ^psi_f[249][7:0];
       end
    500: begin
         out_reg[7:0] <= psi_f[250][15:8];
         parity_reg <= ^psi_f[250][15:8];
       end
    501: begin
         out_reg[7:0] <= psi_f[250][7:0];
         parity_reg <= ^psi_f[250][7:0];
       end
    502: begin
         out_reg[7:0] <= psi_f[251][15:8];
         parity_reg <= ^psi_f[251][15:8];
       end
    503: begin
         out_reg[7:0] <= psi_f[251][7:0];
         parity_reg <= ^psi_f[251][7:0];
       end
    504: begin
         out_reg[7:0] <= psi_f[252][15:8];
         parity_reg <= ^psi_f[252][15:8];
       end
    505: begin
         out_reg[7:0] <= psi_f[252][7:0];
         parity_reg <= ^psi_f[252][7:0];
       end
    506: begin
         out_reg[7:0] <= psi_f[253][15:8];
         parity_reg <= ^psi_f[253][15:8];
       end
    507: begin
         out_reg[7:0] <= psi_f[253][7:0];
         parity_reg <= ^psi_f[253][7:0];
       end
    508: begin
         out_reg[7:0] <= psi_f[254][15:8];
         parity_reg <= ^psi_f[254][15:8];
       end
    509: begin
         out_reg[7:0] <= psi_f[254][7:0];
         parity_reg <= ^psi_f[254][7:0];
       end
    510: begin
         out_reg[7:0] <= psi_f[255][15:8];
         parity_reg <= ^psi_f[255][15:8];
       end
    511: begin
         out_reg[7:0] <= psi_f[255][7:0];
         parity_reg <= ^psi_f[255][7:0];
       end
    512: begin
         out_reg[7:0] <= psi_f[256][15:8];
         parity_reg <= ^psi_f[256][15:8];
       end
    513: begin
         out_reg[7:0] <= psi_f[256][7:0];
         parity_reg <= ^psi_f[256][7:0];
       end
    514: begin
         out_reg[7:0] <= psi_f[257][15:8];
         parity_reg <= ^psi_f[257][15:8];
       end
    515: begin
         out_reg[7:0] <= psi_f[257][7:0];
         parity_reg <= ^psi_f[257][7:0];
       end
    516: begin
         out_reg[7:0] <= psi_f[258][15:8];
         parity_reg <= ^psi_f[258][15:8];
       end
    517: begin
         out_reg[7:0] <= psi_f[258][7:0];
         parity_reg <= ^psi_f[258][7:0];
       end
    518: begin
         out_reg[7:0] <= psi_f[259][15:8];
         parity_reg <= ^psi_f[259][15:8];
       end
    519: begin
         out_reg[7:0] <= psi_f[259][7:0];
         parity_reg <= ^psi_f[259][7:0];
       end
    520: begin
         out_reg[7:0] <= psi_f[260][15:8];
         parity_reg <= ^psi_f[260][15:8];
       end
    521: begin
         out_reg[7:0] <= psi_f[260][7:0];
         parity_reg <= ^psi_f[260][7:0];
       end
    522: begin
         out_reg[7:0] <= psi_f[261][15:8];
         parity_reg <= ^psi_f[261][15:8];
       end
    523: begin
         out_reg[7:0] <= psi_f[261][7:0];
         parity_reg <= ^psi_f[261][7:0];
       end
    524: begin
         out_reg[7:0] <= psi_f[262][15:8];
         parity_reg <= ^psi_f[262][15:8];
       end
    525: begin
         out_reg[7:0] <= psi_f[262][7:0];
         parity_reg <= ^psi_f[262][7:0];
       end
    526: begin
         out_reg[7:0] <= psi_f[263][15:8];
         parity_reg <= ^psi_f[263][15:8];
       end
    527: begin
         out_reg[7:0] <= psi_f[263][7:0];
         parity_reg <= ^psi_f[263][7:0];
       end
    528: begin
         out_reg[7:0] <= psi_f[264][15:8];
         parity_reg <= ^psi_f[264][15:8];
       end
    529: begin
         out_reg[7:0] <= psi_f[264][7:0];
         parity_reg <= ^psi_f[264][7:0];
       end
    530: begin
         out_reg[7:0] <= psi_f[265][15:8];
         parity_reg <= ^psi_f[265][15:8];
       end
    531: begin
         out_reg[7:0] <= psi_f[265][7:0];
         parity_reg <= ^psi_f[265][7:0];
       end
    532: begin
         out_reg[7:0] <= psi_f[266][15:8];
         parity_reg <= ^psi_f[266][15:8];
       end
    533: begin
         out_reg[7:0] <= psi_f[266][7:0];
         parity_reg <= ^psi_f[266][7:0];
       end
    534: begin
         out_reg[7:0] <= psi_f[267][15:8];
         parity_reg <= ^psi_f[267][15:8];
       end
    535: begin
         out_reg[7:0] <= psi_f[267][7:0];
         parity_reg <= ^psi_f[267][7:0];
       end
    536: begin
         out_reg[7:0] <= psi_f[268][15:8];
         parity_reg <= ^psi_f[268][15:8];
       end
    537: begin
         out_reg[7:0] <= psi_f[268][7:0];
         parity_reg <= ^psi_f[268][7:0];
       end
    538: begin
         out_reg[7:0] <= psi_f[269][15:8];
         parity_reg <= ^psi_f[269][15:8];
       end
    539: begin
         out_reg[7:0] <= psi_f[269][7:0];
         parity_reg <= ^psi_f[269][7:0];
       end
    540: begin
         out_reg[7:0] <= psi_f[270][15:8];
         parity_reg <= ^psi_f[270][15:8];
       end
    541: begin
         out_reg[7:0] <= psi_f[270][7:0];
         parity_reg <= ^psi_f[270][7:0];
       end
    542: begin
         out_reg[7:0] <= psi_f[271][15:8];
         parity_reg <= ^psi_f[271][15:8];
       end
    543: begin
         out_reg[7:0] <= psi_f[271][7:0];
         parity_reg <= ^psi_f[271][7:0];
       end
    544: begin
         out_reg[7:0] <= psi_f[272][15:8];
         parity_reg <= ^psi_f[272][15:8];
       end
    545: begin
         out_reg[7:0] <= psi_f[272][7:0];
         parity_reg <= ^psi_f[272][7:0];
       end
    546: begin
         out_reg[7:0] <= psi_f[273][15:8];
         parity_reg <= ^psi_f[273][15:8];
       end
    547: begin
         out_reg[7:0] <= psi_f[273][7:0];
         parity_reg <= ^psi_f[273][7:0];
       end
    548: begin
         out_reg[7:0] <= psi_f[274][15:8];
         parity_reg <= ^psi_f[274][15:8];
       end
    549: begin
         out_reg[7:0] <= psi_f[274][7:0];
         parity_reg <= ^psi_f[274][7:0];
       end
    550: begin
         out_reg[7:0] <= psi_f[275][15:8];
         parity_reg <= ^psi_f[275][15:8];
       end
    551: begin
         out_reg[7:0] <= psi_f[275][7:0];
         parity_reg <= ^psi_f[275][7:0];
       end
    552: begin
         out_reg[7:0] <= psi_f[276][15:8];
         parity_reg <= ^psi_f[276][15:8];
       end
    553: begin
         out_reg[7:0] <= psi_f[276][7:0];
         parity_reg <= ^psi_f[276][7:0];
       end
    554: begin
         out_reg[7:0] <= psi_f[277][15:8];
         parity_reg <= ^psi_f[277][15:8];
       end
    555: begin
         out_reg[7:0] <= psi_f[277][7:0];
         parity_reg <= ^psi_f[277][7:0];
       end
    556: begin
         out_reg[7:0] <= psi_f[278][15:8];
         parity_reg <= ^psi_f[278][15:8];
       end
    557: begin
         out_reg[7:0] <= psi_f[278][7:0];
         parity_reg <= ^psi_f[278][7:0];
       end
    558: begin
         out_reg[7:0] <= psi_f[279][15:8];
         parity_reg <= ^psi_f[279][15:8];
       end
    559: begin
         out_reg[7:0] <= psi_f[279][7:0];
         parity_reg <= ^psi_f[279][7:0];
       end
    560: begin
         out_reg[7:0] <= psi_f[280][15:8];
         parity_reg <= ^psi_f[280][15:8];
       end
    561: begin
         out_reg[7:0] <= psi_f[280][7:0];
         parity_reg <= ^psi_f[280][7:0];
       end
    562: begin
         out_reg[7:0] <= psi_f[281][15:8];
         parity_reg <= ^psi_f[281][15:8];
       end
    563: begin
         out_reg[7:0] <= psi_f[281][7:0];
         parity_reg <= ^psi_f[281][7:0];
       end
    564: begin
         out_reg[7:0] <= psi_f[282][15:8];
         parity_reg <= ^psi_f[282][15:8];
       end
    565: begin
         out_reg[7:0] <= psi_f[282][7:0];
         parity_reg <= ^psi_f[282][7:0];
       end
    566: begin
         out_reg[7:0] <= psi_f[283][15:8];
         parity_reg <= ^psi_f[283][15:8];
       end
    567: begin
         out_reg[7:0] <= psi_f[283][7:0];
         parity_reg <= ^psi_f[283][7:0];
       end
    568: begin
         out_reg[7:0] <= psi_f[284][15:8];
         parity_reg <= ^psi_f[284][15:8];
       end
    569: begin
         out_reg[7:0] <= psi_f[284][7:0];
         parity_reg <= ^psi_f[284][7:0];
       end
    570: begin
         out_reg[7:0] <= psi_f[285][15:8];
         parity_reg <= ^psi_f[285][15:8];
       end
    571: begin
         out_reg[7:0] <= psi_f[285][7:0];
         parity_reg <= ^psi_f[285][7:0];
       end
    572: begin
         out_reg[7:0] <= psi_f[286][15:8];
         parity_reg <= ^psi_f[286][15:8];
       end
    573: begin
         out_reg[7:0] <= psi_f[286][7:0];
         parity_reg <= ^psi_f[286][7:0];
       end
    574: begin
         out_reg[7:0] <= psi_f[287][15:8];
         parity_reg <= ^psi_f[287][15:8];
       end
    575: begin
         out_reg[7:0] <= psi_f[287][7:0];
         parity_reg <= ^psi_f[287][7:0];
       end
    default: out_reg[7:0] <= 8'b00000000;
    endcase
    i_num = i_num + 1;
end
endmodule